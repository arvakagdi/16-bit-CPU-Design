
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Mux is
	Port ( ALUout: IN std_logic_vector (31 downto 0);
	       IRout: IN std_logic_vector (15 downto 0);
	       Sel2: IN std_logic; -- select line for the multiplexer.
	       MuxOut: OUT std_logic_vector(31 downto 0)); -- output the selected input (A for Sel=0) 
end Mux;

architecture behavior of Mux is 
begin

process(ALUout, IRout ,Sel2) 

begin

if (Sel2 = '0') then MuxOut<= ALUout ; 
elsif (Sel2 = '1') then MuxOut<= "0000000000000000" & IRout ; 
end if;

end process;
end behavior;